library verilog;
use verilog.vl_types.all;
entity RISCV_tb is
end RISCV_tb;
